library IEEE;
use IEEE.std_logic_1164.ALL;

entity top is
	port (Clock_50		:	in		std_logic;
			Reset 	:	in		std_logic;
			SW 		:	in		std_logic_vector(9 downto 0);
			LEDR		:	out	std_logic_vector(9 downto 0);
			HEX0		:	out	std_logic_vector(6 downto 0);
			HEX1		:	out	std_logic_vector(6 downto 0);
			HEX2		:	out	std_logic_vector(6 downto 0);
			HEX3		:	out	std_logic_vector(6 downto 0);
			HEX4		:	out	std_logic_vector(6 downto 0);
			HEX5		:	out	std_logic_vector(6 downto 0);
			GPIO_0	:	out	std_logic_vector(15 downto 0);
			KEY		:	in		std_logic_vector(3 downto 0)
			);
end entity;

architecture top_arch of top is

	component char_decoder is
	port (BIN_IN	:	in 	std_logic_vector	(3 downto 0);
			HEX_OUT	:	out 	std_logic_vector	(6 downto 0));
	end component;
	
	component clock_div_prec is
		port (Clock_in		:		in		std_logic;
				Reset 		: 		in		std_logic;
				Sel			: 		in		std_logic_vector (1 downto 0);
				Clock_out	:		out	std_logic);
	end component;

	component computer is
   port  ( clock          : in   std_logic;
				reset          : in   std_logic;
				halted			:	out	std_logic;
				
				port_in_00     : in   std_logic_vector (7 downto 0);
				port_in_01     : in   std_logic_vector (7 downto 0);
				
				port_out_00    : out  std_logic_vector (7 downto 0);
				port_out_01    : out  std_logic_vector (7 downto 0);
				port_out_02    : out  std_logic_vector (7 downto 0);
				port_out_03    : out  std_logic_vector (7 downto 0);
				port_out_04    : out  std_logic_vector (7 downto 0);
				port_out_05    : out  std_logic_vector (7 downto 0);
				
				port_in_02     : in   std_logic_vector (7 downto 0);	
				port_in_03     : in   std_logic_vector (7 downto 0);
				port_in_04     : in   std_logic_vector (7 downto 0);
				port_in_05     : in   std_logic_vector (7 downto 0);
				port_in_06     : in   std_logic_vector (7 downto 0);               
				port_in_07     : in   std_logic_vector (7 downto 0);
				port_in_08     : in   std_logic_vector (7 downto 0);
				port_in_09     : in   std_logic_vector (7 downto 0);
				port_in_10     : in   std_logic_vector (7 downto 0);
				port_in_11     : in   std_logic_vector (7 downto 0);
				port_in_12     : in   std_logic_vector (7 downto 0);
				port_in_13     : in   std_logic_vector (7 downto 0);
				port_in_14     : in   std_logic_vector (7 downto 0);
				port_in_15     : in   std_logic_vector (7 downto 0);                                                                   
				
				port_out_06    : out  std_logic_vector (7 downto 0);
				port_out_07    : out  std_logic_vector (7 downto 0);
				port_out_08    : out  std_logic_vector (7 downto 0);
				port_out_09    : out  std_logic_vector (7 downto 0);
				port_out_10    : out  std_logic_vector (7 downto 0);
				port_out_11    : out  std_logic_vector (7 downto 0);
				port_out_12    : out  std_logic_vector (7 downto 0);
				port_out_13    : out  std_logic_vector (7 downto 0);
				port_out_14    : out  std_logic_vector (7 downto 0);
				port_out_15    : out  std_logic_vector (7 downto 0)
	);
	end component;
	
	signal clock : std_logic;
	
	signal portA,portB,portC,portD,portE	:	std_logic_vector (7 downto 0);
	
	signal nothing1,nothing2,nothing3,nothing4,nothing5,nothing6,nothing7,nothing8,nothing9,nothing10 : std_logic_vector(7 downto 0);
	
	signal halted	: std_logic;
	
begin

	COMP	:	computer port map (	clock,Reset,halted,
											SW(7 downto 0),("0000"&KEY(3 downto 0)),LEDR(7 downto 0),
											portA,portB,portC,portD,portE,
											
											x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
											nothing1,nothing2,nothing3,nothing4,nothing5,nothing6,nothing7,nothing8,nothing9,nothing10
	);

	

	CLOCK_DIV	:	clock_div_prec port map (Clock_50,Reset,SW(9 downto 8),clock);
	
	CHAR_PORTAL	:	char_decoder port map(portA(3 downto 0),HEX0(6 downto 0));
	CHAR_PORTAH :	char_decoder port map(portA(7 downto 4),HEX1(6 downto 0));
	CHAR_PORTBL	:	char_decoder port map(portB(3 downto 0),HEX2(6 downto 0));
	CHAR_PORTBH :	char_decoder port map(portB(7 downto 4),HEX3(6 downto 0));
	CHAR_PORTCL	:	char_decoder port map(portC(3 downto 0),HEX4(6 downto 0));
	CHAR_PORTCH :	char_decoder port map(portC(7 downto 4),HEX5(6 downto 0));
	
	GPIO_0(15 downto 8) <= portE;
	GPIO_0(7 downto 0) <= portD;
	
	LEDR(9) <= halted;
	
end architecture;